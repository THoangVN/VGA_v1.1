module water_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [29:0] color_data
	);

	(* romstyle = "M9K" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		10'b0000000000: color_data = 30'b101001101111011101111111001011;
		10'b0000000001: color_data = 30'b011101011110100111111101100011;
		10'b0000000010: color_data = 30'b011100001110100011111110001011;
		10'b0000000011: color_data = 30'b100000111110111000111110110011;
		10'b0000000100: color_data = 30'b100000001110110010111110110111;
		10'b0000000101: color_data = 30'b011110011110110001111110101011;
		10'b0000000110: color_data = 30'b101100111111011000111111001011;
		10'b0000000111: color_data = 30'b110001001111011111111111010011;
		10'b0000001000: color_data = 30'b011001101110011000111101011111;
		10'b0000001001: color_data = 30'b010101101110000101111100110111;
		10'b0000001010: color_data = 30'b010100111110000100111100100111;
		10'b0000001011: color_data = 30'b010101111110000010111100011111;
		10'b0000001100: color_data = 30'b010101001110000011111100101111;
		10'b0000001101: color_data = 30'b010110111110000001111100101011;
		10'b0000001110: color_data = 30'b010110111110001101111100110011;
		10'b0000001111: color_data = 30'b101100101111011011111111000111;
		10'b0000010000: color_data = 30'b101011011111100011111111101111;
		10'b0000010001: color_data = 30'b011101001110100100111101010011;
		10'b0000010010: color_data = 30'b011100001110100010111101110111;
		10'b0000010011: color_data = 30'b100001001110111000111110101011;
		10'b0000010100: color_data = 30'b011111111110110011111110110011;
		10'b0000010101: color_data = 30'b011110011110110010111110100111;
		10'b0000010110: color_data = 30'b101101011111011001111111001111;
		10'b0000010111: color_data = 30'b101111111111011110111111000011;
		10'b0000011000: color_data = 30'b011010111110011001111101010011;
		10'b0000011001: color_data = 30'b010101111110000011111100110011;
		10'b0000011010: color_data = 30'b010101001110000011111100100111;
		10'b0000011011: color_data = 30'b010101101110000011111100011111;
		10'b0000011100: color_data = 30'b010101001110000101111100101011;
		10'b0000011101: color_data = 30'b010101111110000010111100011111;
		10'b0000011110: color_data = 30'b010101101110001101111100110111;
		10'b0000011111: color_data = 30'b101011111111011000111110111011;

		10'b0000100000: color_data = 30'b100001101110111011111110001111;
		10'b0000100001: color_data = 30'b010011111101111110111100010011;
		10'b0000100010: color_data = 30'b010110111110001100111100111111;
		10'b0000100011: color_data = 30'b011101001110101000111110000111;
		10'b0000100100: color_data = 30'b010111011110001101111100111111;
		10'b0000100101: color_data = 30'b010101101110000111111100100111;
		10'b0000100110: color_data = 30'b011101001110100100111101010011;
		10'b0000100111: color_data = 30'b100010101110111100111101111111;
		10'b0000101000: color_data = 30'b011011011110100001111101110111;
		10'b0000101001: color_data = 30'b011110011110101011111110101011;
		10'b0000101010: color_data = 30'b011010011110011001111101011111;
		10'b0000101011: color_data = 30'b011010011110011100111101110111;
		10'b0000101100: color_data = 30'b011011001110011110111101110111;
		10'b0000101101: color_data = 30'b011011101110011100111101011111;
		10'b0000101110: color_data = 30'b011100011110101000111110100011;
		10'b0000101111: color_data = 30'b100010001111000011111110101111;
		10'b0000110000: color_data = 30'b100001001110111000111101111111;
		10'b0000110001: color_data = 30'b010011101101111111111100001011;
		10'b0000110010: color_data = 30'b010110111110001100111100111011;
		10'b0000110011: color_data = 30'b011101011110100011111101111111;
		10'b0000110100: color_data = 30'b010111111110001011111101001011;
		10'b0000110101: color_data = 30'b010101101110000111111100101011;
		10'b0000110110: color_data = 30'b011110011110100100111101100111;
		10'b0000110111: color_data = 30'b100001111110110111111101111111;
		10'b0000111000: color_data = 30'b011011001110011111111101111011;
		10'b0000111001: color_data = 30'b011101011110101001111110010111;
		10'b0000111010: color_data = 30'b011001101110011010111101010011;
		10'b0000111011: color_data = 30'b011010111110011101111101101011;
		10'b0000111100: color_data = 30'b011010101110011101111101111011;
		10'b0000111101: color_data = 30'b011010111110011101111101101011;
		10'b0000111110: color_data = 30'b011101101110100111111110100111;
		10'b0000111111: color_data = 30'b100001111111000001111110100111;

		10'b0001000000: color_data = 30'b100001111110111001111101111011;
		10'b0001000001: color_data = 30'b010100001101111100111100011111;
		10'b0001000010: color_data = 30'b011010111110011100111101111011;
		10'b0001000011: color_data = 30'b011110101110101100111110011111;
		10'b0001000100: color_data = 30'b010110001110001001111100110011;
		10'b0001000101: color_data = 30'b010101101110000011111100011111;
		10'b0001000110: color_data = 30'b010100011110000001111100100111;
		10'b0001000111: color_data = 30'b100011011110111110111110011011;
		10'b0001001000: color_data = 30'b100010001110101110111101010111;
		10'b0001001001: color_data = 30'b011100111110100011111110001111;
		10'b0001001010: color_data = 30'b100001111110111011111110101111;
		10'b0001001011: color_data = 30'b011110011110110001111110010011;
		10'b0001001100: color_data = 30'b011011111110100011111101111111;
		10'b0001001101: color_data = 30'b011110001110101011111110001011;
		10'b0001001110: color_data = 30'b011010111110011011111101101111;
		10'b0001001111: color_data = 30'b011000001110001110111100101011;
		10'b0001010000: color_data = 30'b011110101110101010111101101111;
		10'b0001010001: color_data = 30'b010011111101111101111100100011;
		10'b0001010010: color_data = 30'b011011001110011101111110000011;
		10'b0001010011: color_data = 30'b011101111110101011111110010111;
		10'b0001010100: color_data = 30'b010110011110001010111100110011;
		10'b0001010101: color_data = 30'b010110111110000010111100110111;
		10'b0001010110: color_data = 30'b010100001110000000111100101011;
		10'b0001010111: color_data = 30'b100100001110111111111110101111;
		10'b0001011000: color_data = 30'b100010011110101011111101100011;
		10'b0001011001: color_data = 30'b011100011110100111111110011111;
		10'b0001011010: color_data = 30'b100001101110111011111110111111;
		10'b0001011011: color_data = 30'b011111001110101101111110011111;
		10'b0001011100: color_data = 30'b011011111110100011111101111111;
		10'b0001011101: color_data = 30'b011110001110101101111110001111;
		10'b0001011110: color_data = 30'b011011001110011001111101110011;
		10'b0001011111: color_data = 30'b010110101110000101111100100111;

		10'b0001100000: color_data = 30'b100101001111001100111110111111;
		10'b0001100001: color_data = 30'b011010011110011101111101100111;
		10'b0001100010: color_data = 30'b011111001110101111111110011011;
		10'b0001100011: color_data = 30'b011101111110100101111110001111;
		10'b0001100100: color_data = 30'b011110011110101010111110010111;
		10'b0001100101: color_data = 30'b011010001110011001111101110011;
		10'b0001100110: color_data = 30'b011010001110011100111101100011;
		10'b0001100111: color_data = 30'b101010011111010101111111000011;
		10'b0001101000: color_data = 30'b101011001111010100111110111011;
		10'b0001101001: color_data = 30'b100010111111000001111110110111;
		10'b0001101010: color_data = 30'b011111111110110110111110111011;
		10'b0001101011: color_data = 30'b010110101110001010111100101011;
		10'b0001101100: color_data = 30'b010011111101111101111100100011;
		10'b0001101101: color_data = 30'b010101111110000101111101000011;
		10'b0001101110: color_data = 30'b011011001110011110111101110111;
		10'b0001101111: color_data = 30'b011100101110100001111101010111;
		10'b0001110000: color_data = 30'b100011101111000010111110101011;
		10'b0001110001: color_data = 30'b011011101110011101111110000111;
		10'b0001110010: color_data = 30'b011110111110101110111110001111;
		10'b0001110011: color_data = 30'b011101011110100110111110000011;
		10'b0001110100: color_data = 30'b011110011110101010111110010111;
		10'b0001110101: color_data = 30'b011010111110010110111101101111;
		10'b0001110110: color_data = 30'b011010001110011100111101100011;
		10'b0001110111: color_data = 30'b101010011111010101111111001011;
		10'b0001111000: color_data = 30'b101011011111010110111110110011;
		10'b0001111001: color_data = 30'b100010001111000011111110110111;
		10'b0001111010: color_data = 30'b100000101110110111111110101111;
		10'b0001111011: color_data = 30'b010110101110001010111100100011;
		10'b0001111100: color_data = 30'b010100011101111111111100101011;
		10'b0001111101: color_data = 30'b010101111110000110111100111011;
		10'b0001111110: color_data = 30'b011010111110100001111110000111;
		10'b0001111111: color_data = 30'b011011111110011110111101011011;

		10'b0010000000: color_data = 30'b100011001111000111111111000111;
		10'b0010000001: color_data = 30'b100000001110110100111111000011;
		10'b0010000010: color_data = 30'b011010111110011001111101011111;
		10'b0010000011: color_data = 30'b010101001110000011111100101111;
		10'b0010000100: color_data = 30'b010110101110000110111100110111;
		10'b0010000101: color_data = 30'b010111011110001110111101000111;
		10'b0010000110: color_data = 30'b100100101111001000111110111011;
		10'b0010000111: color_data = 30'b100010101110111011111110010011;
		10'b0010001000: color_data = 30'b011111001110110100111110011111;
		10'b0010001001: color_data = 30'b100001101110111010111110110011;
		10'b0010001010: color_data = 30'b100100111111000101111110100011;
		10'b0010001011: color_data = 30'b100110001111001010111110101111;
		10'b0010001100: color_data = 30'b011000101110001011111100101111;
		10'b0010001101: color_data = 30'b010111011110001011111100100111;
		10'b0010001110: color_data = 30'b100001111110110111111101110111;
		10'b0010001111: color_data = 30'b101111101111101000111111011011;
		10'b0010010000: color_data = 30'b100100111111001001111110110111;
		10'b0010010001: color_data = 30'b011111101110110100111111000011;
		10'b0010010010: color_data = 30'b011001101110010111111101100111;
		10'b0010010011: color_data = 30'b010101001110000000111100101111;
		10'b0010010100: color_data = 30'b010110011110001000111100110011;
		10'b0010010101: color_data = 30'b010111001110001111111101000111;
		10'b0010010110: color_data = 30'b100101011111001001111111000011;
		10'b0010010111: color_data = 30'b100001011110111010111110001011;
		10'b0010011000: color_data = 30'b011111011110110000111110100111;
		10'b0010011001: color_data = 30'b100001011110111010111110110011;
		10'b0010011010: color_data = 30'b100100001111000110111110101011;
		10'b0010011011: color_data = 30'b100100101111000111111110011111;
		10'b0010011100: color_data = 30'b011000101110001011111100101111;
		10'b0010011101: color_data = 30'b010110101110001011111100110111;
		10'b0010011110: color_data = 30'b100001111110111000111110000011;
		10'b0010011111: color_data = 30'b110000101111100110111111011011;

		10'b0010100000: color_data = 30'b100111101111010100111111011011;
		10'b0010100001: color_data = 30'b011101001110101000111101101011;
		10'b0010100010: color_data = 30'b010101111110000110111100101011;
		10'b0010100011: color_data = 30'b010111101110001000111101000011;
		10'b0010100100: color_data = 30'b010110111110001000111100101111;
		10'b0010100101: color_data = 30'b100011011110111101111110010111;
		10'b0010100110: color_data = 30'b100001101110111101111110010011;
		10'b0010100111: color_data = 30'b010100111110000100111100011111;
		10'b0010101000: color_data = 30'b011101001110100111111110011011;
		10'b0010101001: color_data = 30'b011011111110100110111101111111;
		10'b0010101010: color_data = 30'b010101011110000111111100001011;
		10'b0010101011: color_data = 30'b100101111111000101111110011111;
		10'b0010101100: color_data = 30'b110001111111100111111111011011;
		10'b0010101101: color_data = 30'b101000101111010000111111001011;
		10'b0010101110: color_data = 30'b100110111111010000111111001011;
		10'b0010101111: color_data = 30'b101101101111011011111111010111;
		10'b0010110000: color_data = 30'b101000111111010110111111001111;
		10'b0010110001: color_data = 30'b011011011110100101111101111011;
		10'b0010110010: color_data = 30'b010110011110000101111100110011;
		10'b0010110011: color_data = 30'b010111011110001000111100110111;
		10'b0010110100: color_data = 30'b010110001110001001111100110011;
		10'b0010110101: color_data = 30'b100100101110111110111110001111;
		10'b0010110110: color_data = 30'b100010011110111110111110011011;
		10'b0010110111: color_data = 30'b010101001110000101111100100011;
		10'b0010111000: color_data = 30'b011101111110100111111110010111;
		10'b0010111001: color_data = 30'b011100001110100010111101111111;
		10'b0010111010: color_data = 30'b010101011110000111111100011011;
		10'b0010111011: color_data = 30'b100110011111000111111110100011;
		10'b0010111100: color_data = 30'b110000111111100111111111001111;
		10'b0010111101: color_data = 30'b101000001111010010111111001111;
		10'b0010111110: color_data = 30'b100110111111001101111110111011;
		10'b0010111111: color_data = 30'b101100011111011001111111001011;

		10'b0011000000: color_data = 30'b100101111111001100111110101111;
		10'b0011000001: color_data = 30'b101101001111011110111111011011;
		10'b0011000010: color_data = 30'b101111001111011011111111011111;
		10'b0011000011: color_data = 30'b101100011111011011111111001111;
		10'b0011000100: color_data = 30'b101011101111100001111111011011;
		10'b0011000101: color_data = 30'b110010111111101101111111011111;
		10'b0011000110: color_data = 30'b011111001110100011111101101011;
		10'b0011000111: color_data = 30'b010100001110000001111100110111;
		10'b0011001000: color_data = 30'b011100101110100110111110001011;
		10'b0011001001: color_data = 30'b100000111110111000111110110011;
		10'b0011001010: color_data = 30'b011000011110010010111101010011;
		10'b0011001011: color_data = 30'b010111101110001110111100111011;
		10'b0011001100: color_data = 30'b101010011111010111111111000111;
		10'b0011001101: color_data = 30'b100000001110110100111110010011;
		10'b0011001110: color_data = 30'b010110001110001010111100111111;
		10'b0011001111: color_data = 30'b010110101110001010111100110011;
		10'b0011010000: color_data = 30'b100101001111001001111110100111;
		10'b0011010001: color_data = 30'b101101001111100011111111011111;
		10'b0011010010: color_data = 30'b101111111111011010111111010111;
		10'b0011010011: color_data = 30'b101011111111011101111111010011;
		10'b0011010100: color_data = 30'b101010101111100001111111010111;
		10'b0011010101: color_data = 30'b110011111111101100111111101011;
		10'b0011010110: color_data = 30'b011110011110100100111101100111;
		10'b0011010111: color_data = 30'b010100001110000001111100110111;
		10'b0011011000: color_data = 30'b011100011110101000111110000111;
		10'b0011011001: color_data = 30'b100000001110111010111110101011;
		10'b0011011010: color_data = 30'b011000001110010001111101001111;
		10'b0011011011: color_data = 30'b010111111110001100111100111111;
		10'b0011011100: color_data = 30'b101001001111010010111110110011;
		10'b0011011101: color_data = 30'b100000011110110011111110010011;
		10'b0011011110: color_data = 30'b010110101110001000111101010111;
		10'b0011011111: color_data = 30'b010111111110001100111101000011;

		10'b0011100000: color_data = 30'b010110001110001000111100011011;
		10'b0011100001: color_data = 30'b100110111111000111111110110011;
		10'b0011100010: color_data = 30'b110111001111110010111111111111;
		10'b0011100011: color_data = 30'b101001111111010100111110101111;
		10'b0011100100: color_data = 30'b100010001110110111111110000111;
		10'b0011100101: color_data = 30'b100111011111001010111110011111;
		10'b0011100110: color_data = 30'b100111011111001110111110111011;
		10'b0011100111: color_data = 30'b100001111111000000111110110111;
		10'b0011101000: color_data = 30'b011011011110100001111101110111;
		10'b0011101001: color_data = 30'b011001011110011010111101110011;
		10'b0011101010: color_data = 30'b011110001110101011111110000011;
		10'b0011101011: color_data = 30'b101001001111010011111110111111;
		10'b0011101100: color_data = 30'b100011111111000100111110110011;
		10'b0011101101: color_data = 30'b010110111110001010111100111011;
		10'b0011101110: color_data = 30'b010101111110000001111100100111;
		10'b0011101111: color_data = 30'b010110101110000010111100101011;
		10'b0011110000: color_data = 30'b010111001110001000111100100111;
		10'b0011110001: color_data = 30'b100111011111001010111110100111;
		10'b0011110010: color_data = 30'b110111001111110011111111101111;
		10'b0011110011: color_data = 30'b101010001111010010111110101111;
		10'b0011110100: color_data = 30'b100001111110111000111110000111;
		10'b0011110101: color_data = 30'b100111101111001101111110100111;
		10'b0011110110: color_data = 30'b100110111111001101111110111011;
		10'b0011110111: color_data = 30'b100001111111000001111110111111;
		10'b0011111000: color_data = 30'b011011101110100000111101110111;
		10'b0011111001: color_data = 30'b011010011110011010111101110011;
		10'b0011111010: color_data = 30'b011111001110101001111110000011;
		10'b0011111011: color_data = 30'b101001011111010100111111000011;
		10'b0011111100: color_data = 30'b100011011111000100111110101111;
		10'b0011111101: color_data = 30'b010110111110001011111100110111;
		10'b0011111110: color_data = 30'b010110011110000001111100011011;
		10'b0011111111: color_data = 30'b010110001110000100111100101111;

		10'b0100000000: color_data = 30'b010100101110000000111100110111;
		10'b0100000001: color_data = 30'b011101001110101001111101110111;
		10'b0100000010: color_data = 30'b101001101111011001111111100011;
		10'b0100000011: color_data = 30'b011110101110101101111110001011;
		10'b0100000100: color_data = 30'b011000001110010011111101010011;
		10'b0100000101: color_data = 30'b011100001110100111111101111111;
		10'b0100000110: color_data = 30'b100101111111001000111111000111;
		10'b0100000111: color_data = 30'b100010001110111100111110000111;
		10'b0100001000: color_data = 30'b100001001110101010111101100111;
		10'b0100001001: color_data = 30'b100001111110101100111101011011;
		10'b0100001010: color_data = 30'b011111001110101101111101011011;
		10'b0100001011: color_data = 30'b100111111111000111111110101111;
		10'b0100001100: color_data = 30'b100001001110110111111110110011;
		10'b0100001101: color_data = 30'b010101111110001000111100101111;
		10'b0100001110: color_data = 30'b010110001110000100111100101111;
		10'b0100001111: color_data = 30'b010110101110000100111100111011;
		10'b0100010000: color_data = 30'b010110001101111111111100110011;
		10'b0100010001: color_data = 30'b011110001110101100111101111011;
		10'b0100010010: color_data = 30'b101001011111011000111111001111;
		10'b0100010011: color_data = 30'b011110011110101011111110000011;
		10'b0100010100: color_data = 30'b011000001110010001111101010011;
		10'b0100010101: color_data = 30'b011101001110101000111110000111;
		10'b0100010110: color_data = 30'b100100111111000111111110111111;
		10'b0100010111: color_data = 30'b100010101110111001111110001111;
		10'b0100011000: color_data = 30'b100001101110101101111101100011;
		10'b0100011001: color_data = 30'b100010001110101011111101010111;
		10'b0100011010: color_data = 30'b011111101110101110111101111011;
		10'b0100011011: color_data = 30'b100111011111001010111110100111;
		10'b0100011100: color_data = 30'b100001111110111010111110100111;
		10'b0100011101: color_data = 30'b010111011110001001111101000011;
		10'b0100011110: color_data = 30'b010110001110000010111100101011;
		10'b0100011111: color_data = 30'b010110101110000100111100110011;

		10'b0100100000: color_data = 30'b011110101110110010111110000111;
		10'b0100100001: color_data = 30'b100111111111010010111111000111;
		10'b0100100010: color_data = 30'b100000101110110101111110101011;
		10'b0100100011: color_data = 30'b011111001110110011111110110011;
		10'b0100100100: color_data = 30'b011111111110111001111110011111;
		10'b0100100101: color_data = 30'b100000111110111100111111001111;
		10'b0100100110: color_data = 30'b011011001110011111111101111011;
		10'b0100100111: color_data = 30'b010100001101111111111100010111;
		10'b0100101000: color_data = 30'b101001101111001011111110011011;
		10'b0100101001: color_data = 30'b101101011111011100111110110111;
		10'b0100101010: color_data = 30'b011000011110001101111100110011;
		10'b0100101011: color_data = 30'b010100111110000011111100110111;
		10'b0100101100: color_data = 30'b100000001110110011111110110011;
		10'b0100101101: color_data = 30'b011001111110010111111101010111;
		10'b0100101110: color_data = 30'b010110011110000011111100101111;
		10'b0100101111: color_data = 30'b010101101110000010111100100111;
		10'b0100110000: color_data = 30'b011111111110110001111110001011;
		10'b0100110001: color_data = 30'b100110111111010100111111000111;
		10'b0100110010: color_data = 30'b011111101110110110111110100111;
		10'b0100110011: color_data = 30'b011111111110110011111110110011;
		10'b0100110100: color_data = 30'b100000111110110111111110100111;
		10'b0100110101: color_data = 30'b100010001110111011111111010011;
		10'b0100110110: color_data = 30'b011011001110011110111101101111;
		10'b0100110111: color_data = 30'b010011011101111110111100000111;
		10'b0100111000: color_data = 30'b101010001111001101111110101011;
		10'b0100111001: color_data = 30'b101101101111011100111111001111;
		10'b0100111010: color_data = 30'b010111011110010000111100100111;
		10'b0100111011: color_data = 30'b010101001110000100111100110011;
		10'b0100111100: color_data = 30'b011110001110110100111110100011;
		10'b0100111101: color_data = 30'b011010101110011000111101011011;
		10'b0100111110: color_data = 30'b010110001110000100111100111111;
		10'b0100111111: color_data = 30'b010110011110000101111100110011;

		10'b0101000000: color_data = 30'b110010101111101110111111110011;
		10'b0101000001: color_data = 30'b101000001111000001111110010011;
		10'b0101000010: color_data = 30'b010100101110000010111100110011;
		10'b0101000011: color_data = 30'b010110111110001100111101000111;
		10'b0101000100: color_data = 30'b010110101110001010111101010011;
		10'b0101000101: color_data = 30'b011101001110100110111110010111;
		10'b0101000110: color_data = 30'b011111101110110010111110110011;
		10'b0101000111: color_data = 30'b011001111110011001111101011011;
		10'b0101001000: color_data = 30'b011111011110111001111101111011;
		10'b0101001001: color_data = 30'b011000001110001101111100111011;
		10'b0101001010: color_data = 30'b010101001110000001111100010011;
		10'b0101001011: color_data = 30'b011100101110100101111101110011;
		10'b0101001100: color_data = 30'b100000001110110100111110110111;
		10'b0101001101: color_data = 30'b011111011110110101111110100011;
		10'b0101001110: color_data = 30'b011110101110101111111110001111;
		10'b0101001111: color_data = 30'b100001001110110111111110001011;
		10'b0101010000: color_data = 30'b110010111111101111111111110111;
		10'b0101010001: color_data = 30'b100110111110111101111110000011;
		10'b0101010010: color_data = 30'b010101001110000011111100101111;
		10'b0101010011: color_data = 30'b010110101110001011111101000011;
		10'b0101010100: color_data = 30'b010110101110001001111100111111;
		10'b0101010101: color_data = 30'b011101001110100101111110011111;
		10'b0101010110: color_data = 30'b011111011110110001111110101111;
		10'b0101010111: color_data = 30'b011010001110011000111101100011;
		10'b0101011000: color_data = 30'b100001011110111111111110010111;
		10'b0101011001: color_data = 30'b011000011110010011111101000011;
		10'b0101011010: color_data = 30'b010101001110000000111100100111;
		10'b0101011011: color_data = 30'b011101001110100011111101101111;
		10'b0101011100: color_data = 30'b100000101110110110111110111111;
		10'b0101011101: color_data = 30'b011110111110110100111110101111;
		10'b0101011110: color_data = 30'b011110111110110000111110011011;
		10'b0101011111: color_data = 30'b100001011110111011111101111111;

		10'b0101100000: color_data = 30'b101011001111011011111110111111;
		10'b0101100001: color_data = 30'b101011111111011110111111000011;
		10'b0101100010: color_data = 30'b011011011110100010111101100011;
		10'b0101100011: color_data = 30'b010101001110000000111100100111;
		10'b0101100100: color_data = 30'b010110011110001001111100101111;
		10'b0101100101: color_data = 30'b010110101110001100111100100111;
		10'b0101100110: color_data = 30'b011100101110100101111101111011;
		10'b0101100111: color_data = 30'b100111111111010001111111001011;
		10'b0101101000: color_data = 30'b101111011111100111111111010111;
		10'b0101101001: color_data = 30'b011111111110101110111101110011;
		10'b0101101010: color_data = 30'b011100001110100011111101110011;
		10'b0101101011: color_data = 30'b011101111110101010111110100111;
		10'b0101101100: color_data = 30'b010111001110001101111100111111;
		10'b0101101101: color_data = 30'b010110101110001011111100110111;
		10'b0101101110: color_data = 30'b011111001110110000111110000011;
		10'b0101101111: color_data = 30'b101100001111011110111111010111;
		10'b0101110000: color_data = 30'b101100011111011100111110111111;
		10'b0101110001: color_data = 30'b101011111111011111111111011011;
		10'b0101110010: color_data = 30'b011011001110011111111101010011;
		10'b0101110011: color_data = 30'b010101001101111110111100100011;
		10'b0101110100: color_data = 30'b010110011110001010111100110111;
		10'b0101110101: color_data = 30'b010110111110001100111100111111;
		10'b0101110110: color_data = 30'b011100111110100110111101101111;
		10'b0101110111: color_data = 30'b100110101111001110111111001111;
		10'b0101111000: color_data = 30'b101110111111100101111111010111;
		10'b0101111001: color_data = 30'b100001001110110011111101111111;
		10'b0101111010: color_data = 30'b011100101110100100111101100111;
		10'b0101111011: color_data = 30'b011110001110101001111110010011;
		10'b0101111100: color_data = 30'b010111101110001111111101000111;
		10'b0101111101: color_data = 30'b010101111110001000111100101111;
		10'b0101111110: color_data = 30'b011111111110110011111110001011;
		10'b0101111111: color_data = 30'b101100001111011110111111010111;

		10'b0110000000: color_data = 30'b011011101110100000111101101111;
		10'b0110000001: color_data = 30'b011101011110100111111101101011;
		10'b0110000010: color_data = 30'b101001001111011011111111000011;
		10'b0110000011: color_data = 30'b011111001110110000111101100011;
		10'b0110000100: color_data = 30'b100110001111010000111111000111;
		10'b0110000101: color_data = 30'b100100111111001011111110110011;
		10'b0110000110: color_data = 30'b100100001111000101111110111111;
		10'b0110000111: color_data = 30'b100110001111001010111110101111;
		10'b0110001000: color_data = 30'b101100011111010110111111000111;
		10'b0110001001: color_data = 30'b101010111111100010111111011111;
		10'b0110001010: color_data = 30'b100111001111001101111110110111;
		10'b0110001011: color_data = 30'b010110111110001011111100101111;
		10'b0110001100: color_data = 30'b010101101101111010111100111011;
		10'b0110001101: color_data = 30'b010101011110000001111100110011;
		10'b0110001110: color_data = 30'b100000111110111000111101101011;
		10'b0110001111: color_data = 30'b011100011110100101111101011111;
		10'b0110010000: color_data = 30'b011011011110011010111101111011;
		10'b0110010001: color_data = 30'b011101101110101010111101110011;
		10'b0110010010: color_data = 30'b101001001111011000111111000011;
		10'b0110010011: color_data = 30'b011111111110110000111101100111;
		10'b0110010100: color_data = 30'b100110001111001110111111000011;
		10'b0110010101: color_data = 30'b100101011111001010111110101011;
		10'b0110010110: color_data = 30'b100011101111000011111110111111;
		10'b0110010111: color_data = 30'b100101001111001101111110101111;
		10'b0110011000: color_data = 30'b101011101111010110111110111111;
		10'b0110011001: color_data = 30'b101011101111100001111111011011;
		10'b0110011010: color_data = 30'b100110011111001100111110011111;
		10'b0110011011: color_data = 30'b010111001110001110111100110111;
		10'b0110011100: color_data = 30'b010011101101111110111100101011;
		10'b0110011101: color_data = 30'b010101011110000100111100100011;
		10'b0110011110: color_data = 30'b100001101110111100111110001011;
		10'b0110011111: color_data = 30'b011101111110100101111110000011;

		10'b0110100000: color_data = 30'b011110111110101101111110101011;
		10'b0110100001: color_data = 30'b010100011110000010111100011111;
		10'b0110100010: color_data = 30'b011110011110101110111101100011;
		10'b0110100011: color_data = 30'b100011101111001000111110110111;
		10'b0110100100: color_data = 30'b100000101110111101111110100111;
		10'b0110100101: color_data = 30'b011110001110101011111110010011;
		10'b0110100110: color_data = 30'b010110011110001011111100101011;
		10'b0110100111: color_data = 30'b011000101110010101111101011111;
		10'b0110101000: color_data = 30'b011010001110011100111101100011;
		10'b0110101001: color_data = 30'b100011101111000101111110001111;
		10'b0110101010: color_data = 30'b101111011111101101111111100111;
		10'b0110101011: color_data = 30'b100101001111000110111110100111;
		10'b0110101100: color_data = 30'b011110001110100111111101001111;
		10'b0110101101: color_data = 30'b100101001111000011111101111111;
		10'b0110101110: color_data = 30'b100010011110110110111101111111;
		10'b0110101111: color_data = 30'b010101001110000101111100100011;
		10'b0110110000: color_data = 30'b011101111110101010111110100111;
		10'b0110110001: color_data = 30'b010100101110000100111100001111;
		10'b0110110010: color_data = 30'b100000011110110100111101111111;
		10'b0110110011: color_data = 30'b100100001111001010111111000011;
		10'b0110110100: color_data = 30'b100000101110111000111110011111;
		10'b0110110101: color_data = 30'b011110101110101011111110001111;
		10'b0110110110: color_data = 30'b010101111110001010111100101111;
		10'b0110110111: color_data = 30'b011001011110010110111101100111;
		10'b0110111000: color_data = 30'b011010001110011100111101010111;
		10'b0110111001: color_data = 30'b100100001111000110111110001011;
		10'b0110111010: color_data = 30'b101111011111101101111111101111;
		10'b0110111011: color_data = 30'b100011011111000100111110001111;
		10'b0110111100: color_data = 30'b011101001110100111111101011011;
		10'b0110111101: color_data = 30'b100110001111001001111110011111;
		10'b0110111110: color_data = 30'b100001101110110110111101111011;
		10'b0110111111: color_data = 30'b010100111110000010111100011011;

		10'b0111000000: color_data = 30'b011111111110110011111110110011;
		10'b0111000001: color_data = 30'b010111011110001101111100111111;
		10'b0111000010: color_data = 30'b100100111111000001111110010111;
		10'b0111000011: color_data = 30'b101101001111011110111111010011;
		10'b0111000100: color_data = 30'b011101111110101011111110010111;
		10'b0111000101: color_data = 30'b010101011110000101111100110111;
		10'b0111000110: color_data = 30'b010111011110001111111100111011;
		10'b0111000111: color_data = 30'b011001101110011110111101101111;
		10'b0111001000: color_data = 30'b011100111110100111111101100111;
		10'b0111001001: color_data = 30'b100100101111000101111111000011;
		10'b0111001010: color_data = 30'b011101001110100111111101111011;
		10'b0111001011: color_data = 30'b011110101110110011111110000011;
		10'b0111001100: color_data = 30'b100111101111010100111111011011;
		10'b0111001101: color_data = 30'b101100011111011111111111100111;
		10'b0111001110: color_data = 30'b100111111111010000111111000011;
		10'b0111001111: color_data = 30'b011111111110110101111110010011;
		10'b0111010000: color_data = 30'b100000001110110100111110110111;
		10'b0111010001: color_data = 30'b010111001110001110111100100111;
		10'b0111010010: color_data = 30'b100101011111000011111110010011;
		10'b0111010011: color_data = 30'b101100111111011101111111011011;
		10'b0111010100: color_data = 30'b011110001110101011111110001011;
		10'b0111010101: color_data = 30'b010101101110000110111100111011;
		10'b0111010110: color_data = 30'b010111101110001111111101001011;
		10'b0111010111: color_data = 30'b011001101110011001111101101011;
		10'b0111011000: color_data = 30'b011101101110101010111101110011;
		10'b0111011001: color_data = 30'b100101001111000101111111000011;
		10'b0111011010: color_data = 30'b011101011110100110111101111011;
		10'b0111011011: color_data = 30'b011111001110110001111110001111;
		10'b0111011100: color_data = 30'b100111001111010010111111010011;
		10'b0111011101: color_data = 30'b101011111111011011111111011011;
		10'b0111011110: color_data = 30'b101000011111010010111111001011;
		10'b0111011111: color_data = 30'b011111111110110100111110011011;

		10'b0111100000: color_data = 30'b100111011111010110111111000111;
		10'b0111100001: color_data = 30'b101001011111011110111111001011;
		10'b0111100010: color_data = 30'b101011001111011000111111000111;
		10'b0111100011: color_data = 30'b101100101111001010111110011011;
		10'b0111100100: color_data = 30'b100111001111010001111111000011;
		10'b0111100101: color_data = 30'b100010111111000010111110101111;
		10'b0111100110: color_data = 30'b100101111111000111111110111111;
		10'b0111100111: color_data = 30'b100011111111000100111110110011;
		10'b0111101000: color_data = 30'b011000001110010000111100111011;
		10'b0111101001: color_data = 30'b010110111110000101111100110111;
		10'b0111101010: color_data = 30'b010110111110000011111100100111;
		10'b0111101011: color_data = 30'b010101011110000101111100110111;
		10'b0111101100: color_data = 30'b011001011110010101111101011111;
		10'b0111101101: color_data = 30'b011100001110100010111110000111;
		10'b0111101110: color_data = 30'b011110101110101101111101110011;
		10'b0111101111: color_data = 30'b101001111111011010111111011111;
		10'b0111110000: color_data = 30'b101000011111011010111111010111;
		10'b0111110001: color_data = 30'b101001011111011011111111001111;
		10'b0111110010: color_data = 30'b101010011111010101111110111011;
		10'b0111110011: color_data = 30'b101100101111001010111110011011;
		10'b0111110100: color_data = 30'b100111011111001110111110111011;
		10'b0111110101: color_data = 30'b100010101111000000111110110011;
		10'b0111110110: color_data = 30'b100100011111001001111110111011;
		10'b0111110111: color_data = 30'b100100011111000101111110110111;
		10'b0111111000: color_data = 30'b011000111110010011111101001111;
		10'b0111111001: color_data = 30'b010110111110000111111101000011;
		10'b0111111010: color_data = 30'b010110011110000100111100100111;
		10'b0111111011: color_data = 30'b010110001110000101111100100111;
		10'b0111111100: color_data = 30'b011001001110010101111101011111;
		10'b0111111101: color_data = 30'b011100001110100010111110000111;
		10'b0111111110: color_data = 30'b011110001110101100111101101111;
		10'b0111111111: color_data = 30'b101001001111011010111111001011;

		10'b1000000000: color_data = 30'b101001011111011111111111011111;
		10'b1000000001: color_data = 30'b011111011110101101111101101111;
		10'b1000000010: color_data = 30'b011011001110100011111101100111;
		10'b1000000011: color_data = 30'b011110011110110000111110100011;
		10'b1000000100: color_data = 30'b100001011110111011111110101011;
		10'b1000000101: color_data = 30'b100001011110111101111110110011;
		10'b1000000110: color_data = 30'b101100111111011011111111010111;
		10'b1000000111: color_data = 30'b101111111111100010111111010111;
		10'b1000001000: color_data = 30'b011001111110011001111101011011;
		10'b1000001001: color_data = 30'b010110001110000010111100101011;
		10'b1000001010: color_data = 30'b010101011110000100111100101011;
		10'b1000001011: color_data = 30'b010110001110000010111100110011;
		10'b1000001100: color_data = 30'b010101111110000001111100101111;
		10'b1000001101: color_data = 30'b010101011110000001111100110011;
		10'b1000001110: color_data = 30'b010110101110001011111100111011;
		10'b1000001111: color_data = 30'b101010101111011001111111001111;
		10'b1000010000: color_data = 30'b101011001111100100111111010111;
		10'b1000010001: color_data = 30'b011111001110101101111101100011;
		10'b1000010010: color_data = 30'b011011011110100000111101100111;
		10'b1000010011: color_data = 30'b011110011110110000111110100011;
		10'b1000010100: color_data = 30'b100001111110111001111110101011;
		10'b1000010101: color_data = 30'b100000011110111101111110111111;
		10'b1000010110: color_data = 30'b101100101111011100111111010011;
		10'b1000010111: color_data = 30'b101111111111100011111111000111;
		10'b1000011000: color_data = 30'b011010001110011010111101010111;
		10'b1000011001: color_data = 30'b010110101110000001111100111011;
		10'b1000011010: color_data = 30'b010110001110000101111100100111;
		10'b1000011011: color_data = 30'b010101111110000100111100100011;
		10'b1000011100: color_data = 30'b010101011110000100111100110011;
		10'b1000011101: color_data = 30'b010110101101111110111100101011;
		10'b1000011110: color_data = 30'b010110001110000111111100110111;
		10'b1000011111: color_data = 30'b101011001111010110111110111011;

		10'b1000100000: color_data = 30'b100011011110111110111110100111;
		10'b1000100001: color_data = 30'b010100011101111101111100100011;
		10'b1000100010: color_data = 30'b010111001110001011111100111111;
		10'b1000100011: color_data = 30'b011101111110100101111110000111;
		10'b1000100100: color_data = 30'b010111111110001011111101010011;
		10'b1000100101: color_data = 30'b010101101110000110111100111011;
		10'b1000100110: color_data = 30'b011101011110100011111101011111;
		10'b1000100111: color_data = 30'b100011001110111100111110001011;
		10'b1000101000: color_data = 30'b011011001110011110111101110111;
		10'b1000101001: color_data = 30'b011110001110101010111110011111;
		10'b1000101010: color_data = 30'b011011101110011100111101101011;
		10'b1000101011: color_data = 30'b011011011110011110111101100011;
		10'b1000101100: color_data = 30'b011100101110011111111110001011;
		10'b1000101101: color_data = 30'b011011011110011111111101110011;
		10'b1000101110: color_data = 30'b011100111110100101111110010011;
		10'b1000101111: color_data = 30'b100011001111000010111110100011;
		10'b1000110000: color_data = 30'b100001111110111100111110010011;
		10'b1000110001: color_data = 30'b010100101101111110111100011111;
		10'b1000110010: color_data = 30'b010111001110001101111101000011;
		10'b1000110011: color_data = 30'b011101001110100101111101111111;
		10'b1000110100: color_data = 30'b010111001110001101111101000011;
		10'b1000110101: color_data = 30'b010110011110000101111100110011;
		10'b1000110110: color_data = 30'b011101111110100101111101011011;
		10'b1000110111: color_data = 30'b100001011110110110111101111011;
		10'b1000111000: color_data = 30'b011010111110011110111101111111;
		10'b1000111001: color_data = 30'b011101001110101000111110001011;
		10'b1000111010: color_data = 30'b011010101110011010111101100011;
		10'b1000111011: color_data = 30'b011011111110011111111101111111;
		10'b1000111100: color_data = 30'b011011101110011111111110000111;
		10'b1000111101: color_data = 30'b011011101110011110111101110011;
		10'b1000111110: color_data = 30'b011011011110101001111101111111;
		10'b1000111111: color_data = 30'b100010011111000001111110011011;

		10'b1001000000: color_data = 30'b100001111110111011111110001011;
		10'b1001000001: color_data = 30'b010011101101111101111100010111;
		10'b1001000010: color_data = 30'b011010001110011001111101110011;
		10'b1001000011: color_data = 30'b011110111110101100111110010011;
		10'b1001000100: color_data = 30'b010101111110001000111100101111;
		10'b1001000101: color_data = 30'b010100111110000001111100110011;
		10'b1001000110: color_data = 30'b010100011110000100111100011011;
		10'b1001000111: color_data = 30'b100011011110111111111110010011;
		10'b1001001000: color_data = 30'b100010001110101111111101100011;
		10'b1001001001: color_data = 30'b011101011110100011111101111111;
		10'b1001001010: color_data = 30'b100001111110111010111111000111;
		10'b1001001011: color_data = 30'b011111101110101100111110011111;
		10'b1001001100: color_data = 30'b011011011110100001111101101011;
		10'b1001001101: color_data = 30'b011110001110101001111110001111;
		10'b1001001110: color_data = 30'b011011001110011100111101110011;
		10'b1001001111: color_data = 30'b010111011110010001111100110111;
		10'b1001010000: color_data = 30'b011101111110101011111101101011;
		10'b1001010001: color_data = 30'b010100101101111110111100100111;
		10'b1001010010: color_data = 30'b011010111110011101111101110011;
		10'b1001010011: color_data = 30'b011101111110101011111110010111;
		10'b1001010100: color_data = 30'b010110111110000111111100111011;
		10'b1001010101: color_data = 30'b010110001110000000111100100011;
		10'b1001010110: color_data = 30'b010100011110000000111100100011;
		10'b1001010111: color_data = 30'b100011011110111110111110011011;
		10'b1001011000: color_data = 30'b100010001110101101111101011111;
		10'b1001011001: color_data = 30'b011100111110100110111101111111;
		10'b1001011010: color_data = 30'b100010001110111011111111010011;
		10'b1001011011: color_data = 30'b011110101110101101111110011011;
		10'b1001011100: color_data = 30'b011011001110100000111101110011;
		10'b1001011101: color_data = 30'b011110011110101100111110001111;
		10'b1001011110: color_data = 30'b011011011110100000111101100111;
		10'b1001011111: color_data = 30'b010101111110000111111100011111;

		10'b1001100000: color_data = 30'b100101101111001100111111000011;
		10'b1001100001: color_data = 30'b011010101110011011111101110111;
		10'b1001100010: color_data = 30'b011111011110110000111110100111;
		10'b1001100011: color_data = 30'b011100101110100110111101111111;
		10'b1001100100: color_data = 30'b011110101110101100111110100111;
		10'b1001100101: color_data = 30'b011010101110011101111101111111;
		10'b1001100110: color_data = 30'b011010111110011111111101101111;
		10'b1001100111: color_data = 30'b101010101111010010111111011011;
		10'b1001101000: color_data = 30'b101011101111010100111110011111;
		10'b1001101001: color_data = 30'b100011011111000001111111000111;
		10'b1001101010: color_data = 30'b100000011110110110111110101011;
		10'b1001101011: color_data = 30'b010111001110001001111100110011;
		10'b1001101100: color_data = 30'b010100101101111101111100101111;
		10'b1001101101: color_data = 30'b010101101110000111111100110011;
		10'b1001101110: color_data = 30'b011011001110011100111101110011;
		10'b1001101111: color_data = 30'b011011011110100010111101100011;
		10'b1001110000: color_data = 30'b100011101111000011111110101111;
		10'b1001110001: color_data = 30'b011011011110011101111101110111;
		10'b1001110010: color_data = 30'b011111001110110001111110011111;
		10'b1001110011: color_data = 30'b011101101110100111111110000111;
		10'b1001110100: color_data = 30'b011101111110101100111110001011;
		10'b1001110101: color_data = 30'b011010111110011010111110000011;
		10'b1001110110: color_data = 30'b011010011110011100111101110111;
		10'b1001110111: color_data = 30'b101010111111010100111111001011;
		10'b1001111000: color_data = 30'b101011011111010011111110101011;
		10'b1001111001: color_data = 30'b100011011111000011111110111111;
		10'b1001111010: color_data = 30'b100000101110110101111110101011;
		10'b1001111011: color_data = 30'b010110011110001001111100100111;
		10'b1001111100: color_data = 30'b010101011101111100111100101111;
		10'b1001111101: color_data = 30'b010101111110000110111100110011;
		10'b1001111110: color_data = 30'b011011111110011100111101110111;
		10'b1001111111: color_data = 30'b011011011110100000111101100111;

		10'b1010000000: color_data = 30'b100010111111000111111110110011;
		10'b1010000001: color_data = 30'b011111001110111000111110111011;
		10'b1010000010: color_data = 30'b011010101110010111111101101111;
		10'b1010000011: color_data = 30'b010100111110000011111100101111;
		10'b1010000100: color_data = 30'b010111011110001001111101000011;
		10'b1010000101: color_data = 30'b010111111110010000111101001011;
		10'b1010000110: color_data = 30'b100011011111000101111110101011;
		10'b1010000111: color_data = 30'b100001111110111010111110011111;
		10'b1010001000: color_data = 30'b011111001110110011111110100111;
		10'b1010001001: color_data = 30'b100001101110111100111110101111;
		10'b1010001010: color_data = 30'b100011011111000010111110101011;
		10'b1010001011: color_data = 30'b100101101111001000111110100111;
		10'b1010001100: color_data = 30'b010111101110001011111100111011;
		10'b1010001101: color_data = 30'b010110001110000111111100101111;
		10'b1010001110: color_data = 30'b100010101110110111111110000111;
		10'b1010001111: color_data = 30'b110000111111100100111111011111;
		10'b1010010000: color_data = 30'b100100101111000110111110110111;
		10'b1010010001: color_data = 30'b100000001110110100111110111011;
		10'b1010010010: color_data = 30'b011001111110011001111101011011;
		10'b1010010011: color_data = 30'b010101101101111111111100111011;
		10'b1010010100: color_data = 30'b010111011110001010111100111011;
		10'b1010010101: color_data = 30'b011001011110001101111101001011;
		10'b1010010110: color_data = 30'b100101011111000110111110111111;
		10'b1010010111: color_data = 30'b100001001110111011111110001011;
		10'b1010011000: color_data = 30'b011110101110110010111110110111;
		10'b1010011001: color_data = 30'b100001101110111011111110110111;
		10'b1010011010: color_data = 30'b100011101111000110111110100111;
		10'b1010011011: color_data = 30'b100101001111000110111110011111;
		10'b1010011100: color_data = 30'b010111101110001110111100111011;
		10'b1010011101: color_data = 30'b010101101110000101111100100111;
		10'b1010011110: color_data = 30'b100001011110111001111110000011;
		10'b1010011111: color_data = 30'b110000101111100101111111100011;

		10'b1010100000: color_data = 30'b101001001111010111111111010011;
		10'b1010100001: color_data = 30'b011100111110100111111110000011;
		10'b1010100010: color_data = 30'b010101101110000011111100011111;
		10'b1010100011: color_data = 30'b010110001110000111111100101111;
		10'b1010100100: color_data = 30'b010110011110001000111101000011;
		10'b1010100101: color_data = 30'b100011101110111001111110001111;
		10'b1010100110: color_data = 30'b100010101110111110111110011011;
		10'b1010100111: color_data = 30'b010100111110000010111100011011;
		10'b1010101000: color_data = 30'b011101011110100110111110100111;
		10'b1010101001: color_data = 30'b011011101110100100111110001011;
		10'b1010101010: color_data = 30'b010101111110001001111100010011;
		10'b1010101011: color_data = 30'b100101101111000111111110100011;
		10'b1010101100: color_data = 30'b110001011111100101111111010011;
		10'b1010101101: color_data = 30'b100110111111010001111110110111;
		10'b1010101110: color_data = 30'b100110001111001111111110110111;
		10'b1010101111: color_data = 30'b101100101111011101111110110111;
		10'b1010110000: color_data = 30'b101000001111010110111111001011;
		10'b1010110001: color_data = 30'b011100001110100111111101111111;
		10'b1010110010: color_data = 30'b010110001110000011111100100011;
		10'b1010110011: color_data = 30'b010110011110001000111100110011;
		10'b1010110100: color_data = 30'b010101111110000111111100100111;
		10'b1010110101: color_data = 30'b100010001110111100111110010011;
		10'b1010110110: color_data = 30'b100010111110111010111110010011;
		10'b1010110111: color_data = 30'b010101011110000101111100011111;
		10'b1010111000: color_data = 30'b011101111110100101111110001111;
		10'b1010111001: color_data = 30'b011100001110100010111101111111;
		10'b1010111010: color_data = 30'b010101111110001001111100011011;
		10'b1010111011: color_data = 30'b100110011111000111111110100011;
		10'b1010111100: color_data = 30'b110001011111100010111111001011;
		10'b1010111101: color_data = 30'b100111011111001111111111001011;
		10'b1010111110: color_data = 30'b100101101111001101111110110011;
		10'b1010111111: color_data = 30'b101101011111011010111110110111;

		10'b1011000000: color_data = 30'b100101011111001100111110101011;
		10'b1011000001: color_data = 30'b101101001111011110111111010011;
		10'b1011000010: color_data = 30'b101110101111011000111111000011;
		10'b1011000011: color_data = 30'b101010111111011010111110111011;
		10'b1011000100: color_data = 30'b101010101111011111111111000111;
		10'b1011000101: color_data = 30'b110011111111101100111111101011;
		10'b1011000110: color_data = 30'b011110111110100100111101110011;
		10'b1011000111: color_data = 30'b010100001110000001111100111011;
		10'b1011001000: color_data = 30'b011100111110100111111110001111;
		10'b1011001001: color_data = 30'b100001011110111000111110110111;
		10'b1011001010: color_data = 30'b011000011110010011111101000011;
		10'b1011001011: color_data = 30'b010111111110001100111100111111;
		10'b1011001100: color_data = 30'b101010011111010110111111001111;
		10'b1011001101: color_data = 30'b100001011110110011111110010111;
		10'b1011001110: color_data = 30'b010110011110001010111100111111;
		10'b1011001111: color_data = 30'b010110101110001011111100110111;
		10'b1011010000: color_data = 30'b100100111111001011111110111011;
		10'b1011010001: color_data = 30'b101101011111100000111111001111;
		10'b1011010010: color_data = 30'b101110101111011000111111000011;
		10'b1011010011: color_data = 30'b101011011111011011111111001011;
		10'b1011010100: color_data = 30'b101010111111011101111111010011;
		10'b1011010101: color_data = 30'b110010011111101111111111101011;
		10'b1011010110: color_data = 30'b011110101110100010111110000011;
		10'b1011010111: color_data = 30'b010011111101111110111100111011;
		10'b1011011000: color_data = 30'b011100101110101000111110010011;
		10'b1011011001: color_data = 30'b100001001110111001111110110111;
		10'b1011011010: color_data = 30'b011000101110010011111101100011;
		10'b1011011011: color_data = 30'b010110111110001100111100111011;
		10'b1011011100: color_data = 30'b101010011111010010111110111011;
		10'b1011011101: color_data = 30'b100001001110110011111110100111;
		10'b1011011110: color_data = 30'b010110111110001100111101000111;
		10'b1011011111: color_data = 30'b010111011110001101111100101111;

		10'b1011100000: color_data = 30'b010111011110001000111100110011;
		10'b1011100001: color_data = 30'b100110001111001001111110011111;
		10'b1011100010: color_data = 30'b110111001111110011111111100111;
		10'b1011100011: color_data = 30'b101010101111010001111110111011;
		10'b1011100100: color_data = 30'b100001011110110111111101110011;
		10'b1011100101: color_data = 30'b101000001111001001111110011111;
		10'b1011100110: color_data = 30'b100111011111001111111111000011;
		10'b1011100111: color_data = 30'b100010111110111110111110101111;
		10'b1011101000: color_data = 30'b011010111110011111111101101111;
		10'b1011101001: color_data = 30'b011001001110011010111110000011;
		10'b1011101010: color_data = 30'b011110001110101001111110001111;
		10'b1011101011: color_data = 30'b101001111111001110111110110111;
		10'b1011101100: color_data = 30'b100011001111000100111110100111;
		10'b1011101101: color_data = 30'b010110111110001011111100101111;
		10'b1011101110: color_data = 30'b010101101110000010111100100111;
		10'b1011101111: color_data = 30'b010110001110000010111100101011;
		10'b1011110000: color_data = 30'b010110001110001000111100101011;
		10'b1011110001: color_data = 30'b101000001111001001111110011111;
		10'b1011110010: color_data = 30'b110111011111110101111111111111;
		10'b1011110011: color_data = 30'b101001111111010100111110100111;
		10'b1011110100: color_data = 30'b100000101110110110111101111011;
		10'b1011110101: color_data = 30'b101000011111001011111110010011;
		10'b1011110110: color_data = 30'b100111011111010000111110111111;
		10'b1011110111: color_data = 30'b100010011110111111111110110111;
		10'b1011111000: color_data = 30'b011010101110100000111101110011;
		10'b1011111001: color_data = 30'b011001111110011010111101110011;
		10'b1011111010: color_data = 30'b011110101110101000111110001111;
		10'b1011111011: color_data = 30'b101000111111010001111110101111;
		10'b1011111100: color_data = 30'b100011101111000110111110101111;
		10'b1011111101: color_data = 30'b010110111110001100111101000111;
		10'b1011111110: color_data = 30'b010101111110000001111100100111;
		10'b1011111111: color_data = 30'b010101111110000011111100101011;

		10'b1100000000: color_data = 30'b010101111110000001111100110111;
		10'b1100000001: color_data = 30'b011101111110101100111101100011;
		10'b1100000010: color_data = 30'b101001001111011010111111011011;
		10'b1100000011: color_data = 30'b011110111110101111111110000111;
		10'b1100000100: color_data = 30'b011000111110010100111101011011;
		10'b1100000101: color_data = 30'b011100101110101001111110000111;
		10'b1100000110: color_data = 30'b100100101111000111111110111111;
		10'b1100000111: color_data = 30'b100000011110111000111101111111;
		10'b1100001000: color_data = 30'b100001111110110000111101110011;
		10'b1100001001: color_data = 30'b100011111110110010111101101011;
		10'b1100001010: color_data = 30'b011111101110101110111101110011;
		10'b1100001011: color_data = 30'b100110001111000101111110011011;
		10'b1100001100: color_data = 30'b100001001110111000111110101011;
		10'b1100001101: color_data = 30'b010110011110001010111100110111;
		10'b1100001110: color_data = 30'b010101111110000011111100110011;
		10'b1100001111: color_data = 30'b010111011110000100111100100111;
		10'b1100010000: color_data = 30'b010101001110000000111100100111;
		10'b1100010001: color_data = 30'b011101101110101100111101101111;
		10'b1100010010: color_data = 30'b101001011111011000111111010111;
		10'b1100010011: color_data = 30'b011110001110101101111101111111;
		10'b1100010100: color_data = 30'b011000001110010011111101010111;
		10'b1100010101: color_data = 30'b011101111110101010111110001111;
		10'b1100010110: color_data = 30'b100100001111000111111110111011;
		10'b1100010111: color_data = 30'b100000101110110110111101101111;
		10'b1100011000: color_data = 30'b100000111110110000111101101011;
		10'b1100011001: color_data = 30'b100010101110110100111101110011;
		10'b1100011010: color_data = 30'b011111111110101101111101111011;
		10'b1100011011: color_data = 30'b100111011111000101111110100111;
		10'b1100011100: color_data = 30'b100001101110111000111110101111;
		10'b1100011101: color_data = 30'b010110111110001010111101000011;
		10'b1100011110: color_data = 30'b010110101110000001111100110011;
		10'b1100011111: color_data = 30'b010110011110000110111100101011;

		10'b1100100000: color_data = 30'b011110111110110011111110001011;
		10'b1100100001: color_data = 30'b100110011111010110111111001011;
		10'b1100100010: color_data = 30'b100000101110110111111110100111;
		10'b1100100011: color_data = 30'b011111111110110011111110110111;
		10'b1100100100: color_data = 30'b011111101110111010111110111011;
		10'b1100100101: color_data = 30'b100001001110111101111111010011;
		10'b1100100110: color_data = 30'b011011101110011110111101111011;
		10'b1100100111: color_data = 30'b010100011101111101111100010011;
		10'b1100101000: color_data = 30'b101000111111001010111110100111;
		10'b1100101001: color_data = 30'b101110011111011011111111010011;
		10'b1100101010: color_data = 30'b011000001110010000111101000011;
		10'b1100101011: color_data = 30'b010101011110000100111100110011;
		10'b1100101100: color_data = 30'b011111001110110100111110010111;
		10'b1100101101: color_data = 30'b011010111110010110111101101011;
		10'b1100101110: color_data = 30'b010101101110000101111100100111;
		10'b1100101111: color_data = 30'b010100101110000001111100100111;
		10'b1100110000: color_data = 30'b100000001110110000111110000011;
		10'b1100110001: color_data = 30'b100101101111010011111111001011;
		10'b1100110010: color_data = 30'b100000011110110110111110101011;
		10'b1100110011: color_data = 30'b011111111110110011111110110111;
		10'b1100110100: color_data = 30'b100000001110110111111110110111;
		10'b1100110101: color_data = 30'b100000101110111101111111010111;
		10'b1100110110: color_data = 30'b011010011110011101111101011111;
		10'b1100110111: color_data = 30'b010010101101111011111100000011;
		10'b1100111000: color_data = 30'b101001001111001011111110100011;
		10'b1100111001: color_data = 30'b101100101111011011111110111111;
		10'b1100111010: color_data = 30'b011000001110010000111101000011;
		10'b1100111011: color_data = 30'b010100101110000100111100101111;
		10'b1100111100: color_data = 30'b011110111110110011111110001011;
		10'b1100111101: color_data = 30'b011010001110011010111101011111;
		10'b1100111110: color_data = 30'b010101111110000011111100101011;
		10'b1100111111: color_data = 30'b010101111110000011111100101011;

		10'b1101000000: color_data = 30'b110010001111101100111111101011;
		10'b1101000001: color_data = 30'b101000001111000100111110010011;
		10'b1101000010: color_data = 30'b010101011110000100111100100011;
		10'b1101000011: color_data = 30'b010111001110001101111100111111;
		10'b1101000100: color_data = 30'b010110111110001100111100111011;
		10'b1101000101: color_data = 30'b011101101110100111111110000111;
		10'b1101000110: color_data = 30'b011110101110110001111110100111;
		10'b1101000111: color_data = 30'b011010101110011010111101110011;
		10'b1101001000: color_data = 30'b100001101110111010111110001011;
		10'b1101001001: color_data = 30'b011000111110010001111100110011;
		10'b1101001010: color_data = 30'b010100011110000000111100011011;
		10'b1101001011: color_data = 30'b011011101110100001111101101011;
		10'b1101001100: color_data = 30'b100000111110110110111110111111;
		10'b1101001101: color_data = 30'b011111011110110100111110110011;
		10'b1101001110: color_data = 30'b011101111110101110111110010011;
		10'b1101001111: color_data = 30'b100001001110111001111110010111;
		10'b1101010000: color_data = 30'b110001101111101101111111110011;
		10'b1101010001: color_data = 30'b100111001111000001111101111011;
		10'b1101010010: color_data = 30'b010100111110000100111100100111;
		10'b1101010011: color_data = 30'b010111001110001101111100111111;
		10'b1101010100: color_data = 30'b010111001110001101111100111111;
		10'b1101010101: color_data = 30'b011101001110100110111110010111;
		10'b1101010110: color_data = 30'b011111101110110001111110101011;
		10'b1101010111: color_data = 30'b011010001110011001111101101111;
		10'b1101011000: color_data = 30'b100001011110111111111110011111;
		10'b1101011001: color_data = 30'b011001101110010010111100111111;
		10'b1101011010: color_data = 30'b010100101101111110111100011111;
		10'b1101011011: color_data = 30'b011100011110100010111101110111;
		10'b1101011100: color_data = 30'b100000011110110100111110101111;
		10'b1101011101: color_data = 30'b011111001110110011111110110011;
		10'b1101011110: color_data = 30'b011101111110101111111110001011;
		10'b1101011111: color_data = 30'b100010011110111010111110010111;

		10'b1101100000: color_data = 30'b101100101111010111111111000111;
		10'b1101100001: color_data = 30'b101100011111011110111111010111;
		10'b1101100010: color_data = 30'b011011111110100001111101001011;
		10'b1101100011: color_data = 30'b010100101101111101111100110011;
		10'b1101100100: color_data = 30'b010110011110000110111100011111;
		10'b1101100101: color_data = 30'b010110001110001000111100100011;
		10'b1101100110: color_data = 30'b011011111110100110111101110011;
		10'b1101100111: color_data = 30'b100110111111010011111110111011;
		10'b1101101000: color_data = 30'b110000111111100110111111100111;
		10'b1101101001: color_data = 30'b100001011110110100111101111011;
		10'b1101101010: color_data = 30'b011011111110100011111101110111;
		10'b1101101011: color_data = 30'b011110011110101011111110101011;
		10'b1101101100: color_data = 30'b010111101110001111111101000111;
		10'b1101101101: color_data = 30'b010110101110001011111100110111;
		10'b1101101110: color_data = 30'b011110111110110001111101111111;
		10'b1101101111: color_data = 30'b101011111111011111111111010111;
		10'b1101110000: color_data = 30'b101011111111011101111111010011;
		10'b1101110001: color_data = 30'b101101001111011110111111010011;
		10'b1101110010: color_data = 30'b011100001110011111111101011111;
		10'b1101110011: color_data = 30'b010100111101111010111100011111;
		10'b1101110100: color_data = 30'b010101011110000110111100100111;
		10'b1101110101: color_data = 30'b010101111110001010111100100111;
		10'b1101110110: color_data = 30'b011100101110100111111101110111;
		10'b1101110111: color_data = 30'b100111001111010011111111001011;
		10'b1101111000: color_data = 30'b110000011111101000111111100111;
		10'b1101111001: color_data = 30'b100010001110111000111110000011;
		10'b1101111010: color_data = 30'b011100011110100011111110000011;
		10'b1101111011: color_data = 30'b011110001110101010111110011111;
		10'b1101111100: color_data = 30'b010111101110001111111101000111;
		10'b1101111101: color_data = 30'b010110101110001011111100110111;
		10'b1101111110: color_data = 30'b011111111110110010111101110111;
		10'b1101111111: color_data = 30'b101011011111011101111111000111;

		10'b1110000000: color_data = 30'b011100101110100011111101101111;
		10'b1110000001: color_data = 30'b011101011110100111111101101011;
		10'b1110000010: color_data = 30'b101001001111011010111111001011;
		10'b1110000011: color_data = 30'b100001001110110101111110000011;
		10'b1110000100: color_data = 30'b100110001111001101111110110111;
		10'b1110000101: color_data = 30'b100011111111000011111110101011;
		10'b1110000110: color_data = 30'b100010101110111110111110011011;
		10'b1110000111: color_data = 30'b100101101111000110111110110011;
		10'b1110001000: color_data = 30'b101011101111010101111111010011;
		10'b1110001001: color_data = 30'b101011011111100010111111010011;
		10'b1110001010: color_data = 30'b100111101111010001111111000011;
		10'b1110001011: color_data = 30'b010111001110001100111100111011;
		10'b1110001100: color_data = 30'b010011011101111110111100101011;
		10'b1110001101: color_data = 30'b010101011110000001111100100011;
		10'b1110001110: color_data = 30'b100001111110111011111110000011;
		10'b1110001111: color_data = 30'b011100111110101000111101101011;
		10'b1110010000: color_data = 30'b011010101110011100111101011111;
		10'b1110010001: color_data = 30'b011110001110101000111101100011;
		10'b1110010010: color_data = 30'b101001011111010111111111000011;
		10'b1110010011: color_data = 30'b100001001110110101111101110111;
		10'b1110010100: color_data = 30'b100101101111001011111110110111;
		10'b1110010101: color_data = 30'b100011111111000101111110101111;
		10'b1110010110: color_data = 30'b100010111110111011111110100111;
		10'b1110010111: color_data = 30'b100100101111000110111110101111;
		10'b1110011000: color_data = 30'b101011101111010011111111000011;
		10'b1110011001: color_data = 30'b101011011111100101111111011011;
		10'b1110011010: color_data = 30'b100110011111010001111110110011;
		10'b1110011011: color_data = 30'b010110111110001011111100100111;
		10'b1110011100: color_data = 30'b010011101101111100111100101011;
		10'b1110011101: color_data = 30'b010100111110000010111100011011;
		10'b1110011110: color_data = 30'b100010001110111110111110001011;
		10'b1110011111: color_data = 30'b011101111110101001111101110011;

		10'b1110100000: color_data = 30'b011111001110101110111110100111;
		10'b1110100001: color_data = 30'b010100111101111111111100011011;
		10'b1110100010: color_data = 30'b011111001110101111111101110011;
		10'b1110100011: color_data = 30'b100100101111001010111110111111;
		10'b1110100100: color_data = 30'b100001011110111101111110111011;
		10'b1110100101: color_data = 30'b011110101110101101111110011011;
		10'b1110100110: color_data = 30'b010110001110001011111100110011;
		10'b1110100111: color_data = 30'b011000101110010101111101011111;
		10'b1110101000: color_data = 30'b011010001110011010111101011111;
		10'b1110101001: color_data = 30'b100100111111001010111110100011;
		10'b1110101010: color_data = 30'b101111101111101100111111100111;
		10'b1110101011: color_data = 30'b100101001111001000111110110111;
		10'b1110101100: color_data = 30'b011110011110101111111101110111;
		10'b1110101101: color_data = 30'b100101001111000110111110000111;
		10'b1110101110: color_data = 30'b100001101110110010111101100111;
		10'b1110101111: color_data = 30'b010101011110000100111100100011;
		10'b1110110000: color_data = 30'b011101101110101000111110010111;
		10'b1110110001: color_data = 30'b010101001110000011111100100111;
		10'b1110110010: color_data = 30'b100000001110110011111101111011;
		10'b1110110011: color_data = 30'b100101011111001101111111001011;
		10'b1110110100: color_data = 30'b100001111110111100111111000011;
		10'b1110110101: color_data = 30'b011110101110101011111110010111;
		10'b1110110110: color_data = 30'b010110101110001011111100110111;
		10'b1110110111: color_data = 30'b011000011110010110111101100011;
		10'b1110111000: color_data = 30'b011001111110011101111101100111;
		10'b1110111001: color_data = 30'b100101101111000111111110011111;
		10'b1110111010: color_data = 30'b101111111111101110111111100011;
		10'b1110111011: color_data = 30'b100100011111000101111110110011;
		10'b1110111100: color_data = 30'b011111001110101111111101111011;
		10'b1110111101: color_data = 30'b100111011111000110111110011011;
		10'b1110111110: color_data = 30'b100010011110110100111101111111;
		10'b1110111111: color_data = 30'b010100111110000100111100100111;

		10'b1111000000: color_data = 30'b011111111110110111111110100011;
		10'b1111000001: color_data = 30'b010110011110001101111100011011;
		10'b1111000010: color_data = 30'b100101011111000000111110101011;
		10'b1111000011: color_data = 30'b101101101111011111111111001111;
		10'b1111000100: color_data = 30'b011110001110101100111110010111;
		10'b1111000101: color_data = 30'b010101111110001000111100101111;
		10'b1111000110: color_data = 30'b010111101110001110111101000011;
		10'b1111000111: color_data = 30'b011001111110011101111101101111;
		10'b1111001000: color_data = 30'b011101001110100101111101110111;
		10'b1111001001: color_data = 30'b100100111111000011111111000111;
		10'b1111001010: color_data = 30'b011101101110100111111101111111;
		10'b1111001011: color_data = 30'b100000001110110010111110011111;
		10'b1111001100: color_data = 30'b100111011111010100111111001111;
		10'b1111001101: color_data = 30'b101011001111011001111111011011;
		10'b1111001110: color_data = 30'b100111011111001110111110110011;
		10'b1111001111: color_data = 30'b011111101110110100111110001111;
		10'b1111010000: color_data = 30'b100000001110110101111110101111;
		10'b1111010001: color_data = 30'b010110011110001101111100011111;
		10'b1111010010: color_data = 30'b100101001111000101111110011011;
		10'b1111010011: color_data = 30'b101101111111011100111111011011;
		10'b1111010100: color_data = 30'b011110101110101101111110011011;
		10'b1111010101: color_data = 30'b010101011110000110111100100111;
		10'b1111010110: color_data = 30'b010111001110001111111101000111;
		10'b1111010111: color_data = 30'b011010001110011100111101011011;
		10'b1111011000: color_data = 30'b011101011110101000111101111111;
		10'b1111011001: color_data = 30'b100101001111000101111110110111;
		10'b1111011010: color_data = 30'b011101011110101000111101111111;
		10'b1111011011: color_data = 30'b100000001110110100111110010011;
		10'b1111011100: color_data = 30'b100111101111010011111111001011;
		10'b1111011101: color_data = 30'b101011001111011001111111011011;
		10'b1111011110: color_data = 30'b100111011111010011111110111111;
		10'b1111011111: color_data = 30'b100000001110110110111110010011;

		10'b1111100000: color_data = 30'b100110001111010001111110110011;
		10'b1111100001: color_data = 30'b101000011111010111111111001111;
		10'b1111100010: color_data = 30'b101010011111010011111110110011;
		10'b1111100011: color_data = 30'b101001101111000001111101110011;
		10'b1111100100: color_data = 30'b100111011111010000111110110111;
		10'b1111100101: color_data = 30'b100011001111000001111110100111;
		10'b1111100110: color_data = 30'b100100011111001000111110111111;
		10'b1111100111: color_data = 30'b100011111111000100111111000011;
		10'b1111101000: color_data = 30'b011000101110010100111101001111;
		10'b1111101001: color_data = 30'b010111111110001011111100110011;
		10'b1111101010: color_data = 30'b010101101110000000111100110011;
		10'b1111101011: color_data = 30'b010110011110000101111100111011;
		10'b1111101100: color_data = 30'b011000101110010011111101010111;
		10'b1111101101: color_data = 30'b011010111110011100111101111011;
		10'b1111101110: color_data = 30'b011110011110101101111101110111;
		10'b1111101111: color_data = 30'b101001001111011010111111011011;
		10'b1111110000: color_data = 30'b100110111111010010111111000111;
		10'b1111110001: color_data = 30'b101000011111010111111111001111;
		10'b1111110010: color_data = 30'b101001001111010001111110100011;
		10'b1111110011: color_data = 30'b101000101111000001111101111011;
		10'b1111110100: color_data = 30'b100111011111001110111110111011;
		10'b1111110101: color_data = 30'b100011011111000001111110100111;
		10'b1111110110: color_data = 30'b100100001111000111111111000011;
		10'b1111110111: color_data = 30'b100100011111000110111111000011;
		10'b1111111000: color_data = 30'b011001011110010101111101010111;
		10'b1111111001: color_data = 30'b011000001110001000111100110111;
		10'b1111111010: color_data = 30'b010110001110000010111100101011;
		10'b1111111011: color_data = 30'b010110101110000100111100110011;
		10'b1111111100: color_data = 30'b011000011110010111111101011111;
		10'b1111111101: color_data = 30'b011011011110011101111101111111;
		10'b1111111110: color_data = 30'b011110001110101100111101101111;
		10'b1111111111: color_data = 30'b101001011111011000111111010111;

		default: color_data = 30'b000000000000000000000000000000;
	endcase
endmodule